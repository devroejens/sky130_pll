**.subckt pll_vco vss vdd vtune Ibias
*+ vco_out<0>,vco_out<1>,vco_out<2>,vco_out<3>,vco_out<4>,vco_out<5>,vco_out<6>,vco_out<7> sdn
*.iopin vss
*.iopin vdd
*.iopin vtune
*.iopin Ibias
*.opin vco_out<0>,vco_out<1>,vco_out<2>,vco_out<3>,vco_out<4>,vco_out<5>,vco_out<6>,vco_out<7>
*.iopin sdn
XM0 Ibias Ibias vss vss sky130_fd_pr__nfet_01v8 L=0.3 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
x5<0> phi<0> vss vss vdd vdd net1<7> sky130_fd_sc_hs__inv_1
x5<1> phi<1> vss vss vdd vdd net1<6> sky130_fd_sc_hs__inv_1
x5<2> phi<2> vss vss vdd vdd net1<5> sky130_fd_sc_hs__inv_1
x5<3> phi<3> vss vss vdd vdd net1<4> sky130_fd_sc_hs__inv_1
x5<4> phi<4> vss vss vdd vdd net1<3> sky130_fd_sc_hs__inv_1
x5<5> phi<5> vss vss vdd vdd net1<2> sky130_fd_sc_hs__inv_1
x5<6> phi<6> vss vss vdd vdd net1<1> sky130_fd_sc_hs__inv_1
x5<7> phi<7> vss vss vdd vdd net1<0> sky130_fd_sc_hs__inv_1
x6<0> net1<7> vss vss vdd vdd net2<7> sky130_fd_sc_hs__inv_2
x6<1> net1<6> vss vss vdd vdd net2<6> sky130_fd_sc_hs__inv_2
x6<2> net1<5> vss vss vdd vdd net2<5> sky130_fd_sc_hs__inv_2
x6<3> net1<4> vss vss vdd vdd net2<4> sky130_fd_sc_hs__inv_2
x6<4> net1<3> vss vss vdd vdd net2<3> sky130_fd_sc_hs__inv_2
x6<5> net1<2> vss vss vdd vdd net2<2> sky130_fd_sc_hs__inv_2
x6<6> net1<1> vss vss vdd vdd net2<1> sky130_fd_sc_hs__inv_2
x6<7> net1<0> vss vss vdd vdd net2<0> sky130_fd_sc_hs__inv_2
x7<0> net2<7> vss vss vdd vdd vco_out<0> sky130_fd_sc_hs__inv_4
x7<1> net2<6> vss vss vdd vdd vco_out<1> sky130_fd_sc_hs__inv_4
x7<2> net2<5> vss vss vdd vdd vco_out<2> sky130_fd_sc_hs__inv_4
x7<3> net2<4> vss vss vdd vdd vco_out<3> sky130_fd_sc_hs__inv_4
x7<4> net2<3> vss vss vdd vdd vco_out<4> sky130_fd_sc_hs__inv_4
x7<5> net2<2> vss vss vdd vdd vco_out<5> sky130_fd_sc_hs__inv_4
x7<6> net2<1> vss vss vdd vdd vco_out<6> sky130_fd_sc_hs__inv_4
x7<7> net2<0> vss vss vdd vdd vco_out<7> sky130_fd_sc_hs__inv_4
x1 phi<0> phi<4> phi<7> phi<3> vdd vtune Ibias vss sdn pll_vco_cell
x2 phi<1> phi<5> phi<0> phi<4> vdd vtune Ibias vss sdn pll_vco_cell
x3 phi<2> phi<6> phi<1> phi<5> vdd vtune Ibias vss sdn pll_vco_cell
x4 phi<3> phi<7> phi<2> phi<6> vdd vtune Ibias vss sdn pll_vco_cell
**** begin user architecture code


.control
save i(@m.${path}xm1.msky130_fd_pr__nfet_01v8[id])
save @m.${path}xm1.msky130_fd_pr__nfet_01v8[gm]
save v(@m.${path}xm1.msky130_fd_pr__nfet_01v8[vds])
save v(@m.${path}xm1.msky130_fd_pr__nfet_01v8[vgs])
save v(@m.${path}xm1.msky130_fd_pr__nfet_01v8[vth])
save v(@m.${path}xm1.msky130_fd_pr__nfet_01v8[vdsat])

save i(@m.${path}xm2.msky130_fd_pr__nfet_01v8[id])
save @m.${path}xm2.msky130_fd_pr__nfet_01v8[gm]
save v(@m.${path}xm2.msky130_fd_pr__nfet_01v8[vds])
save v(@m.${path}xm2.msky130_fd_pr__nfet_01v8[vgs])
save v(@m.${path}xm2.msky130_fd_pr__nfet_01v8[vth])
save v(@m.${path}xm2.msky130_fd_pr__nfet_01v8[vdsat])
.endc


**** end user architecture code
**.ends

* expanding   symbol:  pll_vco_cell/xschem/pll_vco_cell.sym # of pins=9
* sym_path: /home/jdv/sky130_pll/pll/pll_vco_cell/xschem/pll_vco_cell.sym
* sch_path: /home/jdv/sky130_pll/pll/pll_vco_cell/xschem/pll_vco_cell.sch
.subckt pll_vco_cell  out_n out_p in_p in_n vdd vtune vbias vss sdn
*.iopin vss
*.iopin vdd
*.ipin in_p
*.ipin in_n
*.iopin vbias
*.opin out_n
*.opin out_p
*.ipin vtune
*.ipin sdn
**** begin user architecture code


*.control
*save i(@m.${path}xm1.msky130_fd_pr__nfet_01v8[id])
*save @m.${path}xm1.msky130_fd_pr__nfet_01v8[gm]
*save v(@m.${path}xm1.msky130_fd_pr__nfet_01v8[vds])
*save v(@m.${path}xm1.msky130_fd_pr__nfet_01v8[vgs])
*save v(@m.${path}xm1.msky130_fd_pr__nfet_01v8[vth])
*save v(@m.${path}xm1.msky130_fd_pr__nfet_01v8[vdsat])

*save i(@m.${path}xm2.msky130_fd_pr__nfet_01v8[id])
*save @m.${path}xm2.msky130_fd_pr__nfet_01v8[gm]
*save v(@m.${path}xm2.msky130_fd_pr__nfet_01v8[vds])
*save v(@m.${path}xm2.msky130_fd_pr__nfet_01v8[vgs])
*save v(@m.${path}xm2.msky130_fd_pr__nfet_01v8[vth])
*save v(@m.${path}xm2.msky130_fd_pr__nfet_01v8[vdsat])
*.endc


**** end user architecture code
XM3 net1 vbias vss vss sky130_fd_pr__nfet_01v8 L=0.3 W=60 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XM10 vbias sdn vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
x1 sdn vss vss vdd vdd net2 sky130_fd_sc_hd__inv_1
x2 sdn vss vss vdd vdd net3 sky130_fd_sc_hd__inv_1
XM4 out_n out_n vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM5 out_p out_p vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM7 out_p out_n vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=16 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM6 out_n out_p vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=16 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM8 out_n net2 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM9 out_p net3 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM1 out_n in_p net1 vss sky130_fd_pr__nfet_01v8 L=0.15 W=16 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM2 out_p in_n net1 vss sky130_fd_pr__nfet_01v8 L=0.15 W=16 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XC1 out_n vtune vss sky130_fd_pr__cap_var_lvt W=7 L=4 VM=3
XC2 out_p vtune vss sky130_fd_pr__cap_var_lvt W=7 L=4 VM=3
.ends

** flattened .save nodes
.end
